module rtc(

);



endmodule
