`timescale 1ns / 1ps

module display(

);

endmodule
