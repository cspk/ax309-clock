`timescale 1ns / 1ps

module clock(
	input wire clk
);

always @ (posedge clk) begin
end

endmodule
