module rtc(
	input sclk,
	input poll_freq,

	output reg ce,

	inout data_io
);



endmodule
