`timescale 1ns / 1ps

module time(

);



endmodule
